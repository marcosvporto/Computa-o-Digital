----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:38:47 03/27/2020 
-- Design Name: 
-- Module Name:    register4 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity register4 is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           D : in  STD_LOGIC_VECTOR(3 downto 0);
           Q : out  STD_LOGIC_VECTOR(3 downto 0)
	 );
end register4;

architecture Behavioral of register4 is

begin

	process (clk)
	begin
		if rising_edge(clk) then
			if (reset = '1') then
				q <= (others => '0');
			else
				Q <= D;
			end if;
		end if;
	end process;

end Behavioral;

